*pmos load inverter

.include /mnt/shared/Docs/Rudra/NITK/sem5/Vlsi_lab/t14y_tsmc_025_level3.txt

mny vndy vy 0 0 cmosn l=1u w=1u
mnx vout vx vndy vndy cmosn l=1u w=1u
mpy vout vy vdd vdd cmosp l = 1u w=1u
mpx vout vx vdd vdd cmosp l = 1u w=1u

v_dd vdd 0 5
v_x vx 0 pulse(0 5 0n 1p 1p 5n 10n)
v_y vy 0 pulse(0 5 2.5n 1p 1p 5n 10n)

cload vout 0 10f

.dc v_x 0 5 0.1
.tran 0.01 40n

.control


.endc
.control
*     foreach x 1u 2u 4u
*     alter m1 w=$x
    run
*     meas tran vmin MIN out FROM=5n to=30n
*     meas tran vmax MAX out FROM=5n to=30n
*     let v10 = vmin  + 0.1*(vmax-vmin)
*     let v90 = vmin  + 0.9*(vmax-vmin)
*     print v10 v90
*
*     meas tran tr TRIG out VAL=v10 RISE=1 TARG out VAL=v90 RISE=1
*     meas tran tf TRIG out VAL=v90 FALL=1 TARG out VAL=v10 FALL=1
*
*     let v_50 = vmin + (vmax-vmin)/2
*
*     meas tran pdhl TRIG vin VAL=2.5 RISE=1 targ out VAL=v_50 FALL=1
*     meas tran pdlh TRIG vin VAL=2.5 FALL=1 TARG out VAL=v_50 RISE=1
*
*     let pd = (pdhl+pdlh)/2
*
*     let slope = deriv(out)
*
*     meas dc voh find out WHEN slope =-1 cross =1
*     meas dc vil find vin WHEN slope = -1 cross = 1
*     meas dc vol find out WHEN slope =-1 cross =2
*     meas dc vih find vin WHEN slope = -1 cross = 2
*
*     let nmh = voh - vih
*     let nml = vil -vol
*     print nmh nml
*     let pwr = (vdd)*(-vdd#branch)
*     meas tran Pavg AVG pwr from=0n to=200n
*     meas tran Pmax MAX pwr from=0n to=200n
*     meas tran Energy INTEG pwr from=0n to=200n
*     end
.endc


.control
    plot tran1.vout vx vy
    plot dc1.vout
.endc
.end
