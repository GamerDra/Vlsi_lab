*NMOS Char

.include /home/rudra/Documents/vlsilab/t14y_tsmc_025_level3.txt
m1 drain gate source bulk cmosn l=1u w=0.5u
vdd drain 0 3.3
vin gate 0 3.3
vss source 0 0
vbb bulk 0 3.3

.dc vin 0 3.3 0.1

.control
foreach vb -2 -1  1 2
alter vbb=$vb
run
end
.endc

.control
foreach iter 1 2 3 4
setplot dc$iter
plot (-vdd#branch)
end
.endc

.end
