*NMOS Characterstics

*includ eth model files
.include /home/vlsilab/UG_students_2025/t14y_tsmc_025_level3.txt

*netist
* m_instance_name drain_mode gate_node
*m` vdd in vaa 0 xmoan l=1u
m1 drain gate 0 0 cmosn l=3u w=20u

vdd drain 0 dc 5
vgg gate 0 dc 5

.dc vgg 0 3.3 0.1 vdd 0 3.3 1


.control
foreach x 1.6e-6 6.4e-6 96e-6
alter m1 l = $x
run
end
.endc

.control
foreach iter 1 2 3
setplot dc$iter
plot -vdd#branch
end
.endc

.control
set filetype=ascii
write output.txt
.endc
.end
